module titulo ( 
	clk,
	set,
	reset,
	j,
	k,
	s,
	r,
	d,
	t,
	selector,
	q,
	qn
	) ;

input  clk;
input  set;
input  reset;
input  j;
input  k;
input  s;
input  r;
input  d;
input  t;
input [1:0] selector;
inout  q;
inout  qn;
