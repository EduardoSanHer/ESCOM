module cr ( 
	clk,
	clr,
	ci,
	cd,
	e,
	ctr,
	q
	) ;

input  clk;
input  clr;
input  ci;
input  cd;
input [6:0] e;
input [2:0] ctr;
inout [6:0] q;
