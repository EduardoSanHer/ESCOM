LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX IS
	PORT(	A,B: IN STD_LOGIC;
			S: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			Z: IN STD_LOGIC
	);
END ENTITY;
ARCHITECTURE A_MUX OF MUX IS
BEGIN
	PROCESS(S)
	BEGIN
		CASE S IS
			WHEN "000" => Z<= A OR B;
			WHEN "001" => Z<= A AND B;
			WHEN "010" => Z<= A NOR B;
			WHEN "011" => Z<= A NAND B;
			WHEN "100" => Z<= A XOR B;
			WHEN "101" => Z<= A XNOR B;
			WHEN "110" => Z<= NOT A;
			WHEN OTHERS => Z<= NOT B;
		END CASE;
	END PROCESS;
	--WITH S SELECT
	--Z <= A OR BS WHEN "000",
		 --A AND B WHEN "001",
		 --A NOR B WHEN "010",
		 --A NAND B WHEN "011",
		 --A XOR B WHEN "100",
		 --A XNOR B WHEN "101",
		 --NOT A WHEN "110",
		 --NOT B WHEN OTHERS;
END A_MUX;
