module ds ( 
	clk,
	x,
	display,
	z
	) ;

input  clk;
input  x;
inout [6:0] display;
inout  z;
