LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PRAC1 IS

	PORT (A,B: IN STD_LOGIC;
		C,D,E,F,G,H,I,J: OUT STD_LOGIC;
		);
END ENTITY;

ARCHITECTURE A_PRAC1 OF PRAC1 IS

BEGIN

	C<= A OR B;
	D<= A AND B;
	E<= A NOR B;
	F<= A NAND B;
	G<= A XOR B;
	H<= A XNOR B;
	I<= NOT A;
	J<= NOT B;

END A_PRAC1;