LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
ENTITY  CUADRO IS
    PORT(A,B,C,D,SEL,REF: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
        DISPLAY: OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
        );
END ENTITY;
ARCHITECTURE A_CUADRO OF CUADRO IS
    SIGNAL DATO: STD_LOGIC_VECTOR (1 DOWNTO 0);
    SIGNAL MA,ME,I: STD_LOGIC;
    BEGIN
    WITH SEL SELECT
    DATO <= A WHEN "00",
            B WHEN "01",
            C WHEN "10",
            D WHEN OTHERS;

    MA <= '1' WHEN (DATO>REF) ELSE '0';
    ME <= '1' WHEN (DATO<REF) ELSE '0';
    I <= '1' WHEN (DATO=REF) ELSE '0';

    DISPLAY <= "0000111" WHEN (MA='1') ELSE
               "0110001" WHEN (ME='1') ELSE
               "0110111";
END A_CUADRO;