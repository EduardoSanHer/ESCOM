module comp ( 
	a,
	b,
	i,
	ma,
	me
	) ;

input [3:0] a;
input [3:0] b;
inout  i;
inout  ma;
inout  me;
