module cod ( 
	i,
	q
	) ;

input [9:0] i;
input [3:0] q;
