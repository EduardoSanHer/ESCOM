module mux ( 
	a,
	b,
	s,
	z
	) ;

input  a;
input  b;
input [2:0] s;
input  z;
