LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMP IS
	PORT(	A,B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			I,MA,ME: OUT STD_LOGIC
	);
END ENTITY;
ARCHITECTURE A_COMP OF COMP IS
BEGIN
	PROCESS(A,B)
		BEGIN
			MA<='0';
			ME<='0';
			I<='0';

			IF(A=B) THEN I<='1';
			ELSIF(A<B) THEN ME<='1';
			ELSE	MA<='1';
			END IF;
		END PROCESS;
END A_COMP;
