module pi ( 
	clk,
	clr,
	ctr,
	e,
	s
	) ;

input  clk;
input  clr;
input  ctr;
input [7:0] e;
inout [7:0] s;
